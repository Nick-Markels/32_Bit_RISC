// -----------------------------------------------------------
//	Module:		32-1 MUX Testbench
//	Author:		Jude Gabriel
//	Contact:	gabriel23@up.edu
//	Date:		March 1, 2022
// ----------------------------------------------------------


`timescale 1ns/1ns

module mux32_to_1_tb;

wire [31:0] z;

reg  [31:0] y31;
reg  [31:0] y30;
reg  [31:0] y29;
reg  [31:0] y28;
reg  [31:0] y27;
reg  [31:0] y26;
reg  [31:0] y25;
reg  [31:0] y24;
reg  [31:0] y23;
reg  [31:0] y22;
reg  [31:0] y21;
reg  [31:0] y20;
reg  [31:0] y19;
reg  [31:0] y18;
reg  [31:0] y17;
reg  [31:0] y16;
reg  [31:0] y15;
reg  [31:0] y14;
reg  [31:0] y13;
reg  [31:0] y12;
reg  [31:0] y11;
reg  [31:0] y10;
reg  [31:0] y9;
reg  [31:0] y8;
reg  [31:0] y7;
reg  [31:0] y6;
reg  [31:0] y5;
reg  [31:0] y4;
reg  [31:0] y3;
reg  [31:0] y2;
reg  [31:0] y1;
reg  [31:0] y0;
reg         s4;
reg         s3;
reg         s2;
reg         s1;
reg         s0;

mux32_to_1 mux(z, y31, y30, y29, y28, y27, y26, y25, y24, y23, 
			y22, y21, y20, y19, y18, y17, y16, y15, y14, 
			y13, y12, y11, y10, y9, y8, y7, y6, y5, y4,
			y3, y2, y1, y0, s4, s3, s2, s1, s0);


initial
  begin
	//Select 00000
	#10 s4 = 1'b0; s3 = 1'b0; s2 = 1'b0; s1 = 1'b0; s0 = 1'b0;
		#10 y31 = 32'h00000000; y30 = 32'h00000000; y29 = 32'h00000000; y28 = 32'h00000000; y27 = 32'h00000000; y26 = 32'h00000000; 
	            y25 = 32'h00000000; y24 = 32'h00000000; y23 = 32'h00000000; y22 = 32'h00000000; y21 = 32'h00000000; y20 = 32'h00000000;
		    y19 = 32'h00000000; y18 = 32'h00000000; y17 = 32'h00000000; y16 = 32'h00000000; y15 = 32'h00000000; y14 = 32'h00000000;
	            y13 = 32'h00000000; y12 = 32'h00000000; y11 = 32'h00000000; y10 = 32'h00000000; y9 = 32'h00000000;  y8 = 32'h00000000;
		    y7 = 32'h00000000;  y6 = 32'h00000000;  y5 = 32'h00000000;  y4 = 32'h00000000;  y3 = 32'h00000000;  y2 = 32'h00000000;
		    y1 = 32'h00000000;  y0 = 32'h00000000;

		#10 y31 = 32'h00000000; y30 = 32'h00000000; y29 = 32'h00000000; y28 = 32'h00000000; y27 = 32'h00000000; y26 = 32'h00000000; 
	            y25 = 32'h00000000; y24 = 32'h00000000; y23 = 32'h00000000; y22 = 32'h00000000; y21 = 32'h00000000; y20 = 32'h00000000;
		    y19 = 32'h00000000; y18 = 32'h00000000; y17 = 32'h00000000; y16 = 32'h00000000; y15 = 32'h00000000; y14 = 32'h00000000;
	            y13 = 32'h00000000; y12 = 32'h00000000; y11 = 32'h00000000; y10 = 32'h00000000; y9 = 32'h00000000;  y8 = 32'h00000000;
		    y7 = 32'h00000000;  y6 = 32'h00000000;  y5 = 32'h00000000;  y4 = 32'h00000000;  y3 = 32'h00000000;  y2 = 32'h00000000;
		    y1 = 32'h00000000;  y0 = 32'hFFFFFFFF;
		
	//Select 00001
	#10 s4 = 1'b0; s3 = 1'b0; s2 = 1'b0; s1 = 1'b0; s0 = 1'b1;
		#10 y31 = 32'h00000000; y30 = 32'h00000000; y29 = 32'h00000000; y28 = 32'h00000000; y27 = 32'h00000000; y26 = 32'h00000000; 
	            y25 = 32'h00000000; y24 = 32'h00000000; y23 = 32'h00000000; y22 = 32'h00000000; y21 = 32'h00000000; y20 = 32'h00000000;
		    y19 = 32'h00000000; y18 = 32'h00000000; y17 = 32'h00000000; y16 = 32'h00000000; y15 = 32'h00000000; y14 = 32'h00000000;
	            y13 = 32'h00000000; y12 = 32'h00000000; y11 = 32'h00000000; y10 = 32'h00000000; y9 = 32'h00000000;  y8 = 32'h00000000;
		    y7 = 32'h00000000;  y6 = 32'h00000000;  y5 = 32'h00000000;  y4 = 32'h00000000;  y3 = 32'h00000000;  y2 = 32'h00000000;
		    y1 = 32'h00000000;  y0 = 32'h00000000;

		#10 y31 = 32'h00000000; y30 = 32'h00000000; y29 = 32'h00000000; y28 = 32'h00000000; y27 = 32'h00000000; y26 = 32'h00000000; 
	            y25 = 32'h00000000; y24 = 32'h00000000; y23 = 32'h00000000; y22 = 32'h00000000; y21 = 32'h00000000; y20 = 32'h00000000;
		    y19 = 32'h00000000; y18 = 32'h00000000; y17 = 32'h00000000; y16 = 32'h00000000; y15 = 32'h00000000; y14 = 32'h00000000;
	            y13 = 32'h00000000; y12 = 32'h00000000; y11 = 32'h00000000; y10 = 32'h00000000; y9 = 32'h00000000;  y8 = 32'h00000000;
		    y7 = 32'h00000000;  y6 = 32'h00000000;  y5 = 32'h00000000;  y4 = 32'h00000000;  y3 = 32'h00000000;  y2 = 32'h00000000;
		    y1 = 32'hFFFFFFFF;  y0 = 32'h00000000;

	//Select 00010
	#10 s4 = 1'b0; s3 = 1'b0; s2 = 1'b0; s1 = 1'b1; s0 = 1'b0;
		#10 y31 = 32'h00000000; y30 = 32'h00000000; y29 = 32'h00000000; y28 = 32'h00000000; y27 = 32'h00000000; y26 = 32'h00000000; 
	            y25 = 32'h00000000; y24 = 32'h00000000; y23 = 32'h00000000; y22 = 32'h00000000; y21 = 32'h00000000; y20 = 32'h00000000;
		    y19 = 32'h00000000; y18 = 32'h00000000; y17 = 32'h00000000; y16 = 32'h00000000; y15 = 32'h00000000; y14 = 32'h00000000;
	            y13 = 32'h00000000; y12 = 32'h00000000; y11 = 32'h00000000; y10 = 32'h00000000; y9 = 32'h00000000;  y8 = 32'h00000000;
		    y7 = 32'h00000000;  y6 = 32'h00000000;  y5 = 32'h00000000;  y4 = 32'h00000000;  y3 = 32'h00000000;  y2 = 32'h00000000;
		    y1 = 32'h00000000;  y0 = 32'h00000000;

		#10 y31 = 32'h00000000; y30 = 32'h00000000; y29 = 32'h00000000; y28 = 32'h00000000; y27 = 32'h00000000; y26 = 32'h00000000; 
	            y25 = 32'h00000000; y24 = 32'h00000000; y23 = 32'h00000000; y22 = 32'h00000000; y21 = 32'h00000000; y20 = 32'h00000000;
		    y19 = 32'h00000000; y18 = 32'h00000000; y17 = 32'h00000000; y16 = 32'h00000000; y15 = 32'h00000000; y14 = 32'h00000000;
	            y13 = 32'h00000000; y12 = 32'h00000000; y11 = 32'h00000000; y10 = 32'h00000000; y9 = 32'h00000000;  y8 = 32'h00000000;
		    y7 = 32'h00000000;  y6 = 32'h00000000;  y5 = 32'h00000000;  y4 = 32'h00000000;  y3 = 32'h00000000;  y2 = 32'hFFFFFFFF;
		    y1 = 32'h00000000;  y0 = 32'h00000000;

	//Select 00011
	#10 s4 = 1'b0; s3 = 1'b0; s2 = 1'b0; s1 = 1'b1; s0 = 1'b1;
		#10 y31 = 32'h00000000; y30 = 32'h00000000; y29 = 32'h00000000; y28 = 32'h00000000; y27 = 32'h00000000; y26 = 32'h00000000; 
	            y25 = 32'h00000000; y24 = 32'h00000000; y23 = 32'h00000000; y22 = 32'h00000000; y21 = 32'h00000000; y20 = 32'h00000000;
		    y19 = 32'h00000000; y18 = 32'h00000000; y17 = 32'h00000000; y16 = 32'h00000000; y15 = 32'h00000000; y14 = 32'h00000000;
	            y13 = 32'h00000000; y12 = 32'h00000000; y11 = 32'h00000000; y10 = 32'h00000000; y9 = 32'h00000000;  y8 = 32'h00000000;
		    y7 = 32'h00000000;  y6 = 32'h00000000;  y5 = 32'h00000000;  y4 = 32'h00000000;  y3 = 32'h00000000;  y2 = 32'h00000000;
		    y1 = 32'h00000000;  y0 = 32'h00000000;

		#10 y31 = 32'h00000000; y30 = 32'h00000000; y29 = 32'h00000000; y28 = 32'h00000000; y27 = 32'h00000000; y26 = 32'h00000000; 
	            y25 = 32'h00000000; y24 = 32'h00000000; y23 = 32'h00000000; y22 = 32'h00000000; y21 = 32'h00000000; y20 = 32'h00000000;
		    y19 = 32'h00000000; y18 = 32'h00000000; y17 = 32'h00000000; y16 = 32'h00000000; y15 = 32'h00000000; y14 = 32'h00000000;
	            y13 = 32'h00000000; y12 = 32'h00000000; y11 = 32'h00000000; y10 = 32'h00000000; y9 = 32'h00000000;  y8 = 32'h00000000;
		    y7 = 32'h00000000;  y6 = 32'h00000000;  y5 = 32'h00000000;  y4 = 32'h00000000;  y3 = 32'hFFFFFFFF;  y2 = 32'h00000000;
		    y1 = 32'h00000000;  y0 = 32'h00000000;


	//Select 00100
	#10 s4 = 1'b0; s3 = 1'b0; s2 = 1'b1; s1 = 1'b0; s0 = 1'b0;
		#10 y31 = 32'h00000000; y30 = 32'h00000000; y29 = 32'h00000000; y28 = 32'h00000000; y27 = 32'h00000000; y26 = 32'h00000000; 
	            y25 = 32'h00000000; y24 = 32'h00000000; y23 = 32'h00000000; y22 = 32'h00000000; y21 = 32'h00000000; y20 = 32'h00000000;
		    y19 = 32'h00000000; y18 = 32'h00000000; y17 = 32'h00000000; y16 = 32'h00000000; y15 = 32'h00000000; y14 = 32'h00000000;
	            y13 = 32'h00000000; y12 = 32'h00000000; y11 = 32'h00000000; y10 = 32'h00000000; y9 = 32'h00000000;  y8 = 32'h00000000;
		    y7 = 32'h00000000;  y6 = 32'h00000000;  y5 = 32'h00000000;  y4 = 32'h00000000;  y3 = 32'h00000000;  y2 = 32'h00000000;
		    y1 = 32'h00000000;  y0 = 32'h00000000;

		#10 y31 = 32'h00000000; y30 = 32'h00000000; y29 = 32'h00000000; y28 = 32'h00000000; y27 = 32'h00000000; y26 = 32'h00000000; 
	            y25 = 32'h00000000; y24 = 32'h00000000; y23 = 32'h00000000; y22 = 32'h00000000; y21 = 32'h00000000; y20 = 32'h00000000;
		    y19 = 32'h00000000; y18 = 32'h00000000; y17 = 32'h00000000; y16 = 32'h00000000; y15 = 32'h00000000; y14 = 32'h00000000;
	            y13 = 32'h00000000; y12 = 32'h00000000; y11 = 32'h00000000; y10 = 32'h00000000; y9 = 32'h00000000;  y8 = 32'h00000000;
		    y7 = 32'h00000000;  y6 = 32'h00000000;  y5 = 32'h00000000;  y4 = 32'hFFFFFFFF;  y3 = 32'h00000000;  y2 = 32'h00000000;
		    y1 = 32'h00000000;  y0 = 32'h00000000;


	//Select 00101
	#10 s4 = 1'b0; s3 = 1'b0; s2 = 1'b1; s1 = 1'b0; s0 = 1'b1;
		#10 y31 = 32'h00000000; y30 = 32'h00000000; y29 = 32'h00000000; y28 = 32'h00000000; y27 = 32'h00000000; y26 = 32'h00000000; 
	            y25 = 32'h00000000; y24 = 32'h00000000; y23 = 32'h00000000; y22 = 32'h00000000; y21 = 32'h00000000; y20 = 32'h00000000;
		    y19 = 32'h00000000; y18 = 32'h00000000; y17 = 32'h00000000; y16 = 32'h00000000; y15 = 32'h00000000; y14 = 32'h00000000;
	            y13 = 32'h00000000; y12 = 32'h00000000; y11 = 32'h00000000; y10 = 32'h00000000; y9 = 32'h00000000;  y8 = 32'h00000000;
		    y7 = 32'h00000000;  y6 = 32'h00000000;  y5 = 32'h00000000;  y4 = 32'h00000000;  y3 = 32'h00000000;  y2 = 32'h00000000;
		    y1 = 32'h00000000;  y0 = 32'h00000000;

		#10 y31 = 32'h00000000; y30 = 32'h00000000; y29 = 32'h00000000; y28 = 32'h00000000; y27 = 32'h00000000; y26 = 32'h00000000; 
	            y25 = 32'h00000000; y24 = 32'h00000000; y23 = 32'h00000000; y22 = 32'h00000000; y21 = 32'h00000000; y20 = 32'h00000000;
		    y19 = 32'h00000000; y18 = 32'h00000000; y17 = 32'h00000000; y16 = 32'h00000000; y15 = 32'h00000000; y14 = 32'h00000000;
	            y13 = 32'h00000000; y12 = 32'h00000000; y11 = 32'h00000000; y10 = 32'h00000000; y9 = 32'h00000000;  y8 = 32'h00000000;
		    y7 = 32'h00000000;  y6 = 32'h00000000;  y5 = 32'hFFFFFFFF;  y4 = 32'h00000000;  y3 = 32'h00000000;  y2 = 32'h00000000;
		    y1 = 32'h00000000;  y0 = 32'h00000000;


	//Select 00110
	#10 s4 = 1'b0; s3 = 1'b0; s2 = 1'b1; s1 = 1'b1; s0 = 1'b0;
		#10 y31 = 32'h00000000; y30 = 32'h00000000; y29 = 32'h00000000; y28 = 32'h00000000; y27 = 32'h00000000; y26 = 32'h00000000; 
	            y25 = 32'h00000000; y24 = 32'h00000000; y23 = 32'h00000000; y22 = 32'h00000000; y21 = 32'h00000000; y20 = 32'h00000000;
		    y19 = 32'h00000000; y18 = 32'h00000000; y17 = 32'h00000000; y16 = 32'h00000000; y15 = 32'h00000000; y14 = 32'h00000000;
	            y13 = 32'h00000000; y12 = 32'h00000000; y11 = 32'h00000000; y10 = 32'h00000000; y9 = 32'h00000000;  y8 = 32'h00000000;
		    y7 = 32'h00000000;  y6 = 32'h00000000;  y5 = 32'h00000000;  y4 = 32'h00000000;  y3 = 32'h00000000;  y2 = 32'h00000000;
		    y1 = 32'h00000000;  y0 = 32'h00000000;

		#10 y31 = 32'h00000000; y30 = 32'h00000000; y29 = 32'h00000000; y28 = 32'h00000000; y27 = 32'h00000000; y26 = 32'h00000000; 
	            y25 = 32'h00000000; y24 = 32'h00000000; y23 = 32'h00000000; y22 = 32'h00000000; y21 = 32'h00000000; y20 = 32'h00000000;
		    y19 = 32'h00000000; y18 = 32'h00000000; y17 = 32'h00000000; y16 = 32'h00000000; y15 = 32'h00000000; y14 = 32'h00000000;
	            y13 = 32'h00000000; y12 = 32'h00000000; y11 = 32'h00000000; y10 = 32'h00000000; y9 = 32'h00000000;  y8 = 32'h00000000;
		    y7 = 32'h00000000;  y6 = 32'hFFFFFFFF;  y5 = 32'h00000000;  y4 = 32'h00000000;  y3 = 32'h00000000;  y2 = 32'h00000000;
		    y1 = 32'h00000000;  y0 = 32'h00000000;	


	//Select 00111
	#10 s4 = 1'b0; s3 = 1'b0; s2 = 1'b1; s1 = 1'b1; s0 = 1'b1;
		#10 y31 = 32'h00000000; y30 = 32'h00000000; y29 = 32'h00000000; y28 = 32'h00000000; y27 = 32'h00000000; y26 = 32'h00000000; 
	            y25 = 32'h00000000; y24 = 32'h00000000; y23 = 32'h00000000; y22 = 32'h00000000; y21 = 32'h00000000; y20 = 32'h00000000;
		    y19 = 32'h00000000; y18 = 32'h00000000; y17 = 32'h00000000; y16 = 32'h00000000; y15 = 32'h00000000; y14 = 32'h00000000;
	            y13 = 32'h00000000; y12 = 32'h00000000; y11 = 32'h00000000; y10 = 32'h00000000; y9 = 32'h00000000;  y8 = 32'h00000000;
		    y7 = 32'h00000000;  y6 = 32'h00000000;  y5 = 32'h00000000;  y4 = 32'h00000000;  y3 = 32'h00000000;  y2 = 32'h00000000;
		    y1 = 32'h00000000;  y0 = 32'h00000000;

		#10 y31 = 32'h00000000; y30 = 32'h00000000; y29 = 32'h00000000; y28 = 32'h00000000; y27 = 32'h00000000; y26 = 32'h00000000; 
	            y25 = 32'h00000000; y24 = 32'h00000000; y23 = 32'h00000000; y22 = 32'h00000000; y21 = 32'h00000000; y20 = 32'h00000000;
		    y19 = 32'h00000000; y18 = 32'h00000000; y17 = 32'h00000000; y16 = 32'h00000000; y15 = 32'h00000000; y14 = 32'h00000000;
	            y13 = 32'h00000000; y12 = 32'h00000000; y11 = 32'h00000000; y10 = 32'h00000000; y9 = 32'h00000000;  y8 = 32'h00000000;
		    y7 = 32'hFFFFFFFF;  y6 = 32'h00000000;  y5 = 32'h00000000;  y4 = 32'h00000000;  y3 = 32'h00000000;  y2 = 32'h00000000;
		    y1 = 32'h00000000;  y0 = 32'h00000000;


	//Select 01000
	#10 s4 = 1'b0; s3 = 1'b1; s2 = 1'b0; s1 = 1'b0; s0 = 1'b0;
		#10 y31 = 32'h00000000; y30 = 32'h00000000; y29 = 32'h00000000; y28 = 32'h00000000; y27 = 32'h00000000; y26 = 32'h00000000; 
	            y25 = 32'h00000000; y24 = 32'h00000000; y23 = 32'h00000000; y22 = 32'h00000000; y21 = 32'h00000000; y20 = 32'h00000000;
		    y19 = 32'h00000000; y18 = 32'h00000000; y17 = 32'h00000000; y16 = 32'h00000000; y15 = 32'h00000000; y14 = 32'h00000000;
	            y13 = 32'h00000000; y12 = 32'h00000000; y11 = 32'h00000000; y10 = 32'h00000000; y9 = 32'h00000000;  y8 = 32'h00000000;
		    y7 = 32'h00000000;  y6 = 32'h00000000;  y5 = 32'h00000000;  y4 = 32'h00000000;  y3 = 32'h00000000;  y2 = 32'h00000000;
		    y1 = 32'h00000000;  y0 = 32'h00000000;

		#10 y31 = 32'h00000000; y30 = 32'h00000000; y29 = 32'h00000000; y28 = 32'h00000000; y27 = 32'h00000000; y26 = 32'h00000000; 
	            y25 = 32'h00000000; y24 = 32'h00000000; y23 = 32'h00000000; y22 = 32'h00000000; y21 = 32'h00000000; y20 = 32'h00000000;
		    y19 = 32'h00000000; y18 = 32'h00000000; y17 = 32'h00000000; y16 = 32'h00000000; y15 = 32'h00000000; y14 = 32'h00000000;
	            y13 = 32'h00000000; y12 = 32'h00000000; y11 = 32'h00000000; y10 = 32'h00000000; y9 = 32'h00000000;  y8 = 32'hFFFFFFFF;
		    y7 = 32'h00000000;  y6 = 32'h00000000;  y5 = 32'h00000000;  y4 = 32'h00000000;  y3 = 32'h00000000;  y2 = 32'h00000000;
		    y1 = 32'h00000000;  y0 = 32'h00000000;


	//Select 01001
	#10 s4 = 1'b0; s3 = 1'b1; s2 = 1'b0; s1 = 1'b0; s0 = 1'b1;
		#10 y31 = 32'h00000000; y30 = 32'h00000000; y29 = 32'h00000000; y28 = 32'h00000000; y27 = 32'h00000000; y26 = 32'h00000000; 
	            y25 = 32'h00000000; y24 = 32'h00000000; y23 = 32'h00000000; y22 = 32'h00000000; y21 = 32'h00000000; y20 = 32'h00000000;
		    y19 = 32'h00000000; y18 = 32'h00000000; y17 = 32'h00000000; y16 = 32'h00000000; y15 = 32'h00000000; y14 = 32'h00000000;
	            y13 = 32'h00000000; y12 = 32'h00000000; y11 = 32'h00000000; y10 = 32'h00000000; y9 = 32'h00000000;  y8 = 32'h00000000;
		    y7 = 32'h00000000;  y6 = 32'h00000000;  y5 = 32'h00000000;  y4 = 32'h00000000;  y3 = 32'h00000000;  y2 = 32'h00000000;
		    y1 = 32'h00000000;  y0 = 32'h00000000;

		#10 y31 = 32'h00000000; y30 = 32'h00000000; y29 = 32'h00000000; y28 = 32'h00000000; y27 = 32'h00000000; y26 = 32'h00000000; 
	            y25 = 32'h00000000; y24 = 32'h00000000; y23 = 32'h00000000; y22 = 32'h00000000; y21 = 32'h00000000; y20 = 32'h00000000;
		    y19 = 32'h00000000; y18 = 32'h00000000; y17 = 32'h00000000; y16 = 32'h00000000; y15 = 32'h00000000; y14 = 32'h00000000;
	            y13 = 32'h00000000; y12 = 32'h00000000; y11 = 32'h00000000; y10 = 32'h00000000; y9 = 32'hFFFFFFFF;  y8 = 32'h00000000;
		    y7 = 32'h00000000;  y6 = 32'h00000000;  y5 = 32'h00000000;  y4 = 32'h00000000;  y3 = 32'h00000000;  y2 = 32'h00000000;
		    y1 = 32'h00000000;  y0 = 32'h00000000;

	//Select 01010
	#10 s4 = 1'b0; s3 = 1'b1; s2 = 1'b0; s1 = 1'b1; s0 = 1'b0;
		#10 y31 = 32'h00000000; y30 = 32'h00000000; y29 = 32'h00000000; y28 = 32'h00000000; y27 = 32'h00000000; y26 = 32'h00000000; 
	            y25 = 32'h00000000; y24 = 32'h00000000; y23 = 32'h00000000; y22 = 32'h00000000; y21 = 32'h00000000; y20 = 32'h00000000;
		    y19 = 32'h00000000; y18 = 32'h00000000; y17 = 32'h00000000; y16 = 32'h00000000; y15 = 32'h00000000; y14 = 32'h00000000;
	            y13 = 32'h00000000; y12 = 32'h00000000; y11 = 32'h00000000; y10 = 32'h00000000; y9 = 32'h00000000;  y8 = 32'h00000000;
		    y7 = 32'h00000000;  y6 = 32'h00000000;  y5 = 32'h00000000;  y4 = 32'h00000000;  y3 = 32'h00000000;  y2 = 32'h00000000;
		    y1 = 32'h00000000;  y0 = 32'h00000000;

		#10 y31 = 32'h00000000; y30 = 32'h00000000; y29 = 32'h00000000; y28 = 32'h00000000; y27 = 32'h00000000; y26 = 32'h00000000; 
	            y25 = 32'h00000000; y24 = 32'h00000000; y23 = 32'h00000000; y22 = 32'h00000000; y21 = 32'h00000000; y20 = 32'h00000000;
		    y19 = 32'h00000000; y18 = 32'h00000000; y17 = 32'h00000000; y16 = 32'h00000000; y15 = 32'h00000000; y14 = 32'h00000000;
	            y13 = 32'h00000000; y12 = 32'h00000000; y11 = 32'h00000000; y10 = 32'hFFFFFFFF; y9 = 32'h00000000;  y8 = 32'h00000000;
		    y7 = 32'h00000000;  y6 = 32'h00000000;  y5 = 32'h00000000;  y4 = 32'h00000000;  y3 = 32'h00000000;  y2 = 32'h00000000;
		    y1 = 32'h00000000;  y0 = 32'h00000000;

	//Select 01011
	#10 s4 = 1'b0; s3 = 1'b1; s2 = 1'b0; s1 = 1'b1; s0 = 1'b1;
		#10 y31 = 32'h00000000; y30 = 32'h00000000; y29 = 32'h00000000; y28 = 32'h00000000; y27 = 32'h00000000; y26 = 32'h00000000; 
	            y25 = 32'h00000000; y24 = 32'h00000000; y23 = 32'h00000000; y22 = 32'h00000000; y21 = 32'h00000000; y20 = 32'h00000000;
		    y19 = 32'h00000000; y18 = 32'h00000000; y17 = 32'h00000000; y16 = 32'h00000000; y15 = 32'h00000000; y14 = 32'h00000000;
	            y13 = 32'h00000000; y12 = 32'h00000000; y11 = 32'h00000000; y10 = 32'h00000000; y9 = 32'h00000000;  y8 = 32'h00000000;
		    y7 = 32'h00000000;  y6 = 32'h00000000;  y5 = 32'h00000000;  y4 = 32'h00000000;  y3 = 32'h00000000;  y2 = 32'h00000000;
		    y1 = 32'h00000000;  y0 = 32'h00000000;

		#10 y31 = 32'h00000000; y30 = 32'h00000000; y29 = 32'h00000000; y28 = 32'h00000000; y27 = 32'h00000000; y26 = 32'h00000000; 
	            y25 = 32'h00000000; y24 = 32'h00000000; y23 = 32'h00000000; y22 = 32'h00000000; y21 = 32'h00000000; y20 = 32'h00000000;
		    y19 = 32'h00000000; y18 = 32'h00000000; y17 = 32'h00000000; y16 = 32'h00000000; y15 = 32'h00000000; y14 = 32'h00000000;
	            y13 = 32'h00000000; y12 = 32'h00000000; y11 = 32'hFFFFFFFF; y10 = 32'h00000000; y9 = 32'h00000000;  y8 = 32'h00000000;
		    y7 = 32'h00000000;  y6 = 32'h00000000;  y5 = 32'h00000000;  y4 = 32'h00000000;  y3 = 32'h00000000;  y2 = 32'h00000000;
		    y1 = 32'h00000000;  y0 = 32'h00000000;

	//Select 01100
	#10 s4 = 1'b0; s3 = 1'b1; s2 = 1'b1; s1 = 1'b0; s0 = 1'b0;
		#10 y31 = 32'h00000000; y30 = 32'h00000000; y29 = 32'h00000000; y28 = 32'h00000000; y27 = 32'h00000000; y26 = 32'h00000000; 
	            y25 = 32'h00000000; y24 = 32'h00000000; y23 = 32'h00000000; y22 = 32'h00000000; y21 = 32'h00000000; y20 = 32'h00000000;
		    y19 = 32'h00000000; y18 = 32'h00000000; y17 = 32'h00000000; y16 = 32'h00000000; y15 = 32'h00000000; y14 = 32'h00000000;
	            y13 = 32'h00000000; y12 = 32'h00000000; y11 = 32'h00000000; y10 = 32'h00000000; y9 = 32'h00000000;  y8 = 32'h00000000;
		    y7 = 32'h00000000;  y6 = 32'h00000000;  y5 = 32'h00000000;  y4 = 32'h00000000;  y3 = 32'h00000000;  y2 = 32'h00000000;
		    y1 = 32'h00000000;  y0 = 32'h00000000;

		#10 y31 = 32'h00000000; y30 = 32'h00000000; y29 = 32'h00000000; y28 = 32'h00000000; y27 = 32'h00000000; y26 = 32'h00000000; 
	            y25 = 32'h00000000; y24 = 32'h00000000; y23 = 32'h00000000; y22 = 32'h00000000; y21 = 32'h00000000; y20 = 32'h00000000;
		    y19 = 32'h00000000; y18 = 32'h00000000; y17 = 32'h00000000; y16 = 32'h00000000; y15 = 32'h00000000; y14 = 32'h00000000;
	            y13 = 32'h00000000; y12 = 32'hFFFFFFFF; y11 = 32'h00000000; y10 = 32'h00000000; y9 = 32'h00000000;  y8 = 32'h00000000;
		    y7 = 32'h00000000;  y6 = 32'h00000000;  y5 = 32'h00000000;  y4 = 32'h00000000;  y3 = 32'h00000000;  y2 = 32'h00000000;
		    y1 = 32'h00000000;  y0 = 32'h00000000;

	//Select 01101
	#10 s4 = 1'b0; s3 = 1'b1; s2 = 1'b1; s1 = 1'b0; s0 = 1'b1;
		#10 y31 = 32'h00000000; y30 = 32'h00000000; y29 = 32'h00000000; y28 = 32'h00000000; y27 = 32'h00000000; y26 = 32'h00000000; 
	            y25 = 32'h00000000; y24 = 32'h00000000; y23 = 32'h00000000; y22 = 32'h00000000; y21 = 32'h00000000; y20 = 32'h00000000;
		    y19 = 32'h00000000; y18 = 32'h00000000; y17 = 32'h00000000; y16 = 32'h00000000; y15 = 32'h00000000; y14 = 32'h00000000;
	            y13 = 32'h00000000; y12 = 32'h00000000; y11 = 32'h00000000; y10 = 32'h00000000; y9 = 32'h00000000;  y8 = 32'h00000000;
		    y7 = 32'h00000000;  y6 = 32'h00000000;  y5 = 32'h00000000;  y4 = 32'h00000000;  y3 = 32'h00000000;  y2 = 32'h00000000;
		    y1 = 32'h00000000;  y0 = 32'h00000000;
		
		#10 y31 = 32'h00000000; y30 = 32'h00000000; y29 = 32'h00000000; y28 = 32'h00000000; y27 = 32'h00000000; y26 = 32'h00000000; 
	            y25 = 32'h00000000; y24 = 32'h00000000; y23 = 32'h00000000; y22 = 32'h00000000; y21 = 32'h00000000; y20 = 32'h00000000;
		    y19 = 32'h00000000; y18 = 32'h00000000; y17 = 32'h00000000; y16 = 32'h00000000; y15 = 32'h00000000; y14 = 32'h00000000;
	            y13 = 32'hFFFFFFFF; y12 = 32'h00000000; y11 = 32'h00000000; y10 = 32'h00000000; y9 = 32'h00000000;  y8 = 32'h00000000;
		    y7 = 32'h00000000;  y6 = 32'h00000000;  y5 = 32'h00000000;  y4 = 32'h00000000;  y3 = 32'h00000000;  y2 = 32'h00000000;
		    y1 = 32'h00000000;  y0 = 32'h00000000;

	//Select 01110
	#10 s4 = 1'b0; s3 = 1'b1; s2 = 1'b1; s1 = 1'b1; s0 = 1'b0;
		#10 y31 = 32'h00000000; y30 = 32'h00000000; y29 = 32'h00000000; y28 = 32'h00000000; y27 = 32'h00000000; y26 = 32'h00000000; 
	            y25 = 32'h00000000; y24 = 32'h00000000; y23 = 32'h00000000; y22 = 32'h00000000; y21 = 32'h00000000; y20 = 32'h00000000;
		    y19 = 32'h00000000; y18 = 32'h00000000; y17 = 32'h00000000; y16 = 32'h00000000; y15 = 32'h00000000; y14 = 32'h00000000;
	            y13 = 32'h00000000; y12 = 32'h00000000; y11 = 32'h00000000; y10 = 32'h00000000; y9 = 32'h00000000;  y8 = 32'h00000000;
		    y7 = 32'h00000000;  y6 = 32'h00000000;  y5 = 32'h00000000;  y4 = 32'h00000000;  y3 = 32'h00000000;  y2 = 32'h00000000;
		    y1 = 32'h00000000;  y0 = 32'h00000000;

		#10 y31 = 32'h00000000; y30 = 32'h00000000; y29 = 32'h00000000; y28 = 32'h00000000; y27 = 32'h00000000; y26 = 32'h00000000; 
	            y25 = 32'h00000000; y24 = 32'h00000000; y23 = 32'h00000000; y22 = 32'h00000000; y21 = 32'h00000000; y20 = 32'h00000000;
		    y19 = 32'h00000000; y18 = 32'h00000000; y17 = 32'h00000000; y16 = 32'h00000000; y15 = 32'h00000000; y14 = 32'hFFFFFFFF;
	            y13 = 32'h00000000; y12 = 32'h00000000; y11 = 32'h00000000; y10 = 32'h00000000; y9 = 32'h00000000;  y8 = 32'h00000000;
		    y7 = 32'h00000000;  y6 = 32'h00000000;  y5 = 32'h00000000;  y4 = 32'h00000000;  y3 = 32'h00000000;  y2 = 32'h00000000;
		    y1 = 32'h00000000;  y0 = 32'h00000000;

	//Select 01111
	#10 s4 = 1'b0; s3 = 1'b1; s2 = 1'b1; s1 = 1'b1; s0 = 1'b1;
		#10 y31 = 32'h00000000; y30 = 32'h00000000; y29 = 32'h00000000; y28 = 32'h00000000; y27 = 32'h00000000; y26 = 32'h00000000; 
	            y25 = 32'h00000000; y24 = 32'h00000000; y23 = 32'h00000000; y22 = 32'h00000000; y21 = 32'h00000000; y20 = 32'h00000000;
		    y19 = 32'h00000000; y18 = 32'h00000000; y17 = 32'h00000000; y16 = 32'h00000000; y15 = 32'h00000000; y14 = 32'h00000000;
	            y13 = 32'h00000000; y12 = 32'h00000000; y11 = 32'h00000000; y10 = 32'h00000000; y9 = 32'h00000000;  y8 = 32'h00000000;
		    y7 = 32'h00000000;  y6 = 32'h00000000;  y5 = 32'h00000000;  y4 = 32'h00000000;  y3 = 32'h00000000;  y2 = 32'h00000000;
		    y1 = 32'h00000000;  y0 = 32'h00000000;

		#10 y31 = 32'h00000000; y30 = 32'h00000000; y29 = 32'h00000000; y28 = 32'h00000000; y27 = 32'h00000000; y26 = 32'h00000000; 
	            y25 = 32'h00000000; y24 = 32'h00000000; y23 = 32'h00000000; y22 = 32'h00000000; y21 = 32'h00000000; y20 = 32'h00000000;
		    y19 = 32'h00000000; y18 = 32'h00000000; y17 = 32'h00000000; y16 = 32'h00000000; y15 = 32'hFFFFFFFF; y14 = 32'h00000000;
	            y13 = 32'h00000000; y12 = 32'h00000000; y11 = 32'h00000000; y10 = 32'h00000000; y9 = 32'h00000000;  y8 = 32'h00000000;
		    y7 = 32'h00000000;  y6 = 32'h00000000;  y5 = 32'h00000000;  y4 = 32'h00000000;  y3 = 32'h00000000;  y2 = 32'h00000000;
		    y1 = 32'h00000000;  y0 = 32'h00000000;

	//Select 10000
	#10 s4 = 1'b1; s3 = 1'b0; s2 = 1'b0; s1 = 1'b0; s0 = 1'b0;
		#10 y31 = 32'h00000000; y30 = 32'h00000000; y29 = 32'h00000000; y28 = 32'h00000000; y27 = 32'h00000000; y26 = 32'h00000000; 
	            y25 = 32'h00000000; y24 = 32'h00000000; y23 = 32'h00000000; y22 = 32'h00000000; y21 = 32'h00000000; y20 = 32'h00000000;
		    y19 = 32'h00000000; y18 = 32'h00000000; y17 = 32'h00000000; y16 = 32'h00000000; y15 = 32'h00000000; y14 = 32'h00000000;
	            y13 = 32'h00000000; y12 = 32'h00000000; y11 = 32'h00000000; y10 = 32'h00000000; y9 = 32'h00000000;  y8 = 32'h00000000;
		    y7 = 32'h00000000;  y6 = 32'h00000000;  y5 = 32'h00000000;  y4 = 32'h00000000;  y3 = 32'h00000000;  y2 = 32'h00000000;
		    y1 = 32'h00000000;  y0 = 32'h00000000;

		#10 y31 = 32'h00000000; y30 = 32'h00000000; y29 = 32'h00000000; y28 = 32'h00000000; y27 = 32'h00000000; y26 = 32'h00000000; 
	            y25 = 32'h00000000; y24 = 32'h00000000; y23 = 32'h00000000; y22 = 32'h00000000; y21 = 32'h00000000; y20 = 32'h00000000;
		    y19 = 32'h00000000; y18 = 32'h00000000; y17 = 32'h00000000; y16 = 32'hFFFFFFFF; y15 = 32'h00000000; y14 = 32'h00000000;
	            y13 = 32'h00000000; y12 = 32'h00000000; y11 = 32'h00000000; y10 = 32'h00000000; y9 = 32'h00000000;  y8 = 32'h00000000;
		    y7 = 32'h00000000;  y6 = 32'h00000000;  y5 = 32'h00000000;  y4 = 32'h00000000;  y3 = 32'h00000000;  y2 = 32'h00000000;
		    y1 = 32'h00000000;  y0 = 32'h00000000;


	//Select 10001
	#10 s4 = 1'b1; s3 = 1'b0; s2 = 1'b0; s1 = 1'b0; s0 = 1'b1;
		#10 y31 = 32'h00000000; y30 = 32'h00000000; y29 = 32'h00000000; y28 = 32'h00000000; y27 = 32'h00000000; y26 = 32'h00000000; 
	            y25 = 32'h00000000; y24 = 32'h00000000; y23 = 32'h00000000; y22 = 32'h00000000; y21 = 32'h00000000; y20 = 32'h00000000;
		    y19 = 32'h00000000; y18 = 32'h00000000; y17 = 32'h00000000; y16 = 32'h00000000; y15 = 32'h00000000; y14 = 32'h00000000;
	            y13 = 32'h00000000; y12 = 32'h00000000; y11 = 32'h00000000; y10 = 32'h00000000; y9 = 32'h00000000;  y8 = 32'h00000000;
		    y7 = 32'h00000000;  y6 = 32'h00000000;  y5 = 32'h00000000;  y4 = 32'h00000000;  y3 = 32'h00000000;  y2 = 32'h00000000;
		    y1 = 32'h00000000;  y0 = 32'h00000000;

		#10 y31 = 32'h00000000; y30 = 32'h00000000; y29 = 32'h00000000; y28 = 32'h00000000; y27 = 32'h00000000; y26 = 32'h00000000; 
	            y25 = 32'h00000000; y24 = 32'h00000000; y23 = 32'h00000000; y22 = 32'h00000000; y21 = 32'h00000000; y20 = 32'h00000000;
		    y19 = 32'h00000000; y18 = 32'h00000000; y17 = 32'hFFFFFFFF; y16 = 32'h00000000; y15 = 32'h00000000; y14 = 32'h00000000;
	            y13 = 32'h00000000; y12 = 32'h00000000; y11 = 32'h00000000; y10 = 32'h00000000; y9 = 32'h00000000;  y8 = 32'h00000000;
		    y7 = 32'h00000000;  y6 = 32'h00000000;  y5 = 32'h00000000;  y4 = 32'h00000000;  y3 = 32'h00000000;  y2 = 32'h00000000;
		    y1 = 32'h00000000;  y0 = 32'h00000000;


	//Select 10010
	#10 s4 = 1'b1; s3 = 1'b0; s2 = 1'b0; s1 = 1'b1; s0 = 1'b0;
		#10 y31 = 32'h00000000; y30 = 32'h00000000; y29 = 32'h00000000; y28 = 32'h00000000; y27 = 32'h00000000; y26 = 32'h00000000; 
	            y25 = 32'h00000000; y24 = 32'h00000000; y23 = 32'h00000000; y22 = 32'h00000000; y21 = 32'h00000000; y20 = 32'h00000000;
		    y19 = 32'h00000000; y18 = 32'h00000000; y17 = 32'h00000000; y16 = 32'h00000000; y15 = 32'h00000000; y14 = 32'h00000000;
	            y13 = 32'h00000000; y12 = 32'h00000000; y11 = 32'h00000000; y10 = 32'h00000000; y9 = 32'h00000000;  y8 = 32'h00000000;
		    y7 = 32'h00000000;  y6 = 32'h00000000;  y5 = 32'h00000000;  y4 = 32'h00000000;  y3 = 32'h00000000;  y2 = 32'h00000000;
		    y1 = 32'h00000000;  y0 = 32'h00000000;

		#10 y31 = 32'h00000000; y30 = 32'h00000000; y29 = 32'h00000000; y28 = 32'h00000000; y27 = 32'h00000000; y26 = 32'h00000000; 
	            y25 = 32'h00000000; y24 = 32'h00000000; y23 = 32'h00000000; y22 = 32'h00000000; y21 = 32'h00000000; y20 = 32'h00000000;
		    y19 = 32'h00000000; y18 = 32'hFFFFFFFF; y17 = 32'h00000000; y16 = 32'h00000000; y15 = 32'h00000000; y14 = 32'h00000000;
	            y13 = 32'h00000000; y12 = 32'h00000000; y11 = 32'h00000000; y10 = 32'h00000000; y9 = 32'h00000000;  y8 = 32'h00000000;
		    y7 = 32'h00000000;  y6 = 32'h00000000;  y5 = 32'h00000000;  y4 = 32'h00000000;  y3 = 32'h00000000;  y2 = 32'h00000000;
		    y1 = 32'h00000000;  y0 = 32'h00000000;


	//Select 10011
	#10 s4 = 1'b1; s3 = 1'b0; s2 = 1'b0; s1 = 1'b1; s0 = 1'b1;
		#10 y31 = 32'h00000000; y30 = 32'h00000000; y29 = 32'h00000000; y28 = 32'h00000000; y27 = 32'h00000000; y26 = 32'h00000000; 
	            y25 = 32'h00000000; y24 = 32'h00000000; y23 = 32'h00000000; y22 = 32'h00000000; y21 = 32'h00000000; y20 = 32'h00000000;
		    y19 = 32'h00000000; y18 = 32'h00000000; y17 = 32'h00000000; y16 = 32'h00000000; y15 = 32'h00000000; y14 = 32'h00000000;
	            y13 = 32'h00000000; y12 = 32'h00000000; y11 = 32'h00000000; y10 = 32'h00000000; y9 = 32'h00000000;  y8 = 32'h00000000;
		    y7 = 32'h00000000;  y6 = 32'h00000000;  y5 = 32'h00000000;  y4 = 32'h00000000;  y3 = 32'h00000000;  y2 = 32'h00000000;
		    y1 = 32'h00000000;  y0 = 32'h00000000;

		#10 y31 = 32'h00000000; y30 = 32'h00000000; y29 = 32'h00000000; y28 = 32'h00000000; y27 = 32'h00000000; y26 = 32'h00000000; 
	            y25 = 32'h00000000; y24 = 32'h00000000; y23 = 32'h00000000; y22 = 32'h00000000; y21 = 32'h00000000; y20 = 32'h00000000;
		    y19 = 32'hFFFFFFFF; y18 = 32'h00000000; y17 = 32'h00000000; y16 = 32'h00000000; y15 = 32'h00000000; y14 = 32'h00000000;
	            y13 = 32'h00000000; y12 = 32'h00000000; y11 = 32'h00000000; y10 = 32'h00000000; y9 = 32'h00000000;  y8 = 32'h00000000;
		    y7 = 32'h00000000;  y6 = 32'h00000000;  y5 = 32'h00000000;  y4 = 32'h00000000;  y3 = 32'h00000000;  y2 = 32'h00000000;
		    y1 = 32'h00000000;  y0 = 32'h00000000;


	//Select 10100
	#10 s4 = 1'b1; s3 = 1'b0; s2 = 1'b1; s1 = 1'b0; s0 = 1'b0;
		#10 y31 = 32'h00000000; y30 = 32'h00000000; y29 = 32'h00000000; y28 = 32'h00000000; y27 = 32'h00000000; y26 = 32'h00000000; 
	            y25 = 32'h00000000; y24 = 32'h00000000; y23 = 32'h00000000; y22 = 32'h00000000; y21 = 32'h00000000; y20 = 32'h00000000;
		    y19 = 32'h00000000; y18 = 32'h00000000; y17 = 32'h00000000; y16 = 32'h00000000; y15 = 32'h00000000; y14 = 32'h00000000;
	            y13 = 32'h00000000; y12 = 32'h00000000; y11 = 32'h00000000; y10 = 32'h00000000; y9 = 32'h00000000;  y8 = 32'h00000000;
		    y7 = 32'h00000000;  y6 = 32'h00000000;  y5 = 32'h00000000;  y4 = 32'h00000000;  y3 = 32'h00000000;  y2 = 32'h00000000;
		    y1 = 32'h00000000;  y0 = 32'h00000000;

		#10 y31 = 32'h00000000; y30 = 32'h00000000; y29 = 32'h00000000; y28 = 32'h00000000; y27 = 32'h00000000; y26 = 32'h00000000; 
	            y25 = 32'h00000000; y24 = 32'h00000000; y23 = 32'h00000000; y22 = 32'h00000000; y21 = 32'h00000000; y20 = 32'hFFFFFFFF;
		    y19 = 32'h00000000; y18 = 32'h00000000; y17 = 32'h00000000; y16 = 32'h00000000; y15 = 32'h00000000; y14 = 32'h00000000;
	            y13 = 32'h00000000; y12 = 32'h00000000; y11 = 32'h00000000; y10 = 32'h00000000; y9 = 32'h00000000;  y8 = 32'h00000000;
		    y7 = 32'h00000000;  y6 = 32'h00000000;  y5 = 32'h00000000;  y4 = 32'h00000000;  y3 = 32'h00000000;  y2 = 32'h00000000;
		    y1 = 32'h00000000;  y0 = 32'h00000000;



	//Select 10101
	#10 s4 = 1'b1; s3 = 1'b0; s2 = 1'b1; s1 = 1'b0; s0 = 1'b1;
		#10 y31 = 32'h00000000; y30 = 32'h00000000; y29 = 32'h00000000; y28 = 32'h00000000; y27 = 32'h00000000; y26 = 32'h00000000; 
	            y25 = 32'h00000000; y24 = 32'h00000000; y23 = 32'h00000000; y22 = 32'h00000000; y21 = 32'h00000000; y20 = 32'h00000000;
		    y19 = 32'h00000000; y18 = 32'h00000000; y17 = 32'h00000000; y16 = 32'h00000000; y15 = 32'h00000000; y14 = 32'h00000000;
	            y13 = 32'h00000000; y12 = 32'h00000000; y11 = 32'h00000000; y10 = 32'h00000000; y9 = 32'h00000000;  y8 = 32'h00000000;
		    y7 = 32'h00000000;  y6 = 32'h00000000;  y5 = 32'h00000000;  y4 = 32'h00000000;  y3 = 32'h00000000;  y2 = 32'h00000000;
		    y1 = 32'h00000000;  y0 = 32'h00000000;

		#10 y31 = 32'h00000000; y30 = 32'h00000000; y29 = 32'h00000000; y28 = 32'h00000000; y27 = 32'h00000000; y26 = 32'h00000000; 
	            y25 = 32'h00000000; y24 = 32'h00000000; y23 = 32'h00000000; y22 = 32'h00000000; y21 = 32'hFFFFFFFF; y20 = 32'h00000000;
		    y19 = 32'h00000000; y18 = 32'h00000000; y17 = 32'h00000000; y16 = 32'h00000000; y15 = 32'h00000000; y14 = 32'h00000000;
	            y13 = 32'h00000000; y12 = 32'h00000000; y11 = 32'h00000000; y10 = 32'h00000000; y9 = 32'h00000000;  y8 = 32'h00000000;
		    y7 = 32'h00000000;  y6 = 32'h00000000;  y5 = 32'h00000000;  y4 = 32'h00000000;  y3 = 32'h00000000;  y2 = 32'h00000000;
		    y1 = 32'h00000000;  y0 = 32'h00000000;

	//Select 10110
	#10 s4 = 1'b1; s3 = 1'b0; s2 = 1'b1; s1 = 1'b1; s0 = 1'b0;
		#10 y31 = 32'h00000000; y30 = 32'h00000000; y29 = 32'h00000000; y28 = 32'h00000000; y27 = 32'h00000000; y26 = 32'h00000000; 
	            y25 = 32'h00000000; y24 = 32'h00000000; y23 = 32'h00000000; y22 = 32'h00000000; y21 = 32'h00000000; y20 = 32'h00000000;
		    y19 = 32'h00000000; y18 = 32'h00000000; y17 = 32'h00000000; y16 = 32'h00000000; y15 = 32'h00000000; y14 = 32'h00000000;
	            y13 = 32'h00000000; y12 = 32'h00000000; y11 = 32'h00000000; y10 = 32'h00000000; y9 = 32'h00000000;  y8 = 32'h00000000;
		    y7 = 32'h00000000;  y6 = 32'h00000000;  y5 = 32'h00000000;  y4 = 32'h00000000;  y3 = 32'h00000000;  y2 = 32'h00000000;
		    y1 = 32'h00000000;  y0 = 32'h00000000;
		
		#10 y31 = 32'h00000000; y30 = 32'h00000000; y29 = 32'h00000000; y28 = 32'h00000000; y27 = 32'h00000000; y26 = 32'h00000000; 
	            y25 = 32'h00000000; y24 = 32'h00000000; y23 = 32'h00000000; y22 = 32'hFFFFFFFF; y21 = 32'h00000000; y20 = 32'h00000000;
		    y19 = 32'h00000000; y18 = 32'h00000000; y17 = 32'h00000000; y16 = 32'h00000000; y15 = 32'h00000000; y14 = 32'h00000000;
	            y13 = 32'h00000000; y12 = 32'h00000000; y11 = 32'h00000000; y10 = 32'h00000000; y9 = 32'h00000000;  y8 = 32'h00000000;
		    y7 = 32'h00000000;  y6 = 32'h00000000;  y5 = 32'h00000000;  y4 = 32'h00000000;  y3 = 32'h00000000;  y2 = 32'h00000000;
		    y1 = 32'h00000000;  y0 = 32'h00000000;
	
	//Select 10111
	#10 s4 = 1'b1; s3 = 1'b0; s2 = 1'b1; s1 = 1'b1; s0 = 1'b1;
		#10 y31 = 32'h00000000; y30 = 32'h00000000; y29 = 32'h00000000; y28 = 32'h00000000; y27 = 32'h00000000; y26 = 32'h00000000; 
	            y25 = 32'h00000000; y24 = 32'h00000000; y23 = 32'h00000000; y22 = 32'h00000000; y21 = 32'h00000000; y20 = 32'h00000000;
		    y19 = 32'h00000000; y18 = 32'h00000000; y17 = 32'h00000000; y16 = 32'h00000000; y15 = 32'h00000000; y14 = 32'h00000000;
	            y13 = 32'h00000000; y12 = 32'h00000000; y11 = 32'h00000000; y10 = 32'h00000000; y9 = 32'h00000000;  y8 = 32'h00000000;
		    y7 = 32'h00000000;  y6 = 32'h00000000;  y5 = 32'h00000000;  y4 = 32'h00000000;  y3 = 32'h00000000;  y2 = 32'h00000000;
		    y1 = 32'h00000000;  y0 = 32'h00000000;

		#10 y31 = 32'h00000000; y30 = 32'h00000000; y29 = 32'h00000000; y28 = 32'h00000000; y27 = 32'h00000000; y26 = 32'h00000000; 
	            y25 = 32'h00000000; y24 = 32'h00000000; y23 = 32'hFFFFFFFF; y22 = 32'h00000000; y21 = 32'h00000000; y20 = 32'h00000000;
		    y19 = 32'h00000000; y18 = 32'h00000000; y17 = 32'h00000000; y16 = 32'h00000000; y15 = 32'h00000000; y14 = 32'h00000000;
	            y13 = 32'h00000000; y12 = 32'h00000000; y11 = 32'h00000000; y10 = 32'h00000000; y9 = 32'h00000000;  y8 = 32'h00000000;
		    y7 = 32'h00000000;  y6 = 32'h00000000;  y5 = 32'h00000000;  y4 = 32'h00000000;  y3 = 32'h00000000;  y2 = 32'h00000000;
		    y1 = 32'h00000000;  y0 = 32'h00000000;


	//Select 11000
	#10 s4 = 1'b1; s3 = 1'b1; s2 = 1'b0; s1 = 1'b0; s0 = 1'b0;
		#10 y31 = 32'h00000000; y30 = 32'h00000000; y29 = 32'h00000000; y28 = 32'h00000000; y27 = 32'h00000000; y26 = 32'h00000000; 
	            y25 = 32'h00000000; y24 = 32'h00000000; y23 = 32'h00000000; y22 = 32'h00000000; y21 = 32'h00000000; y20 = 32'h00000000;
		    y19 = 32'h00000000; y18 = 32'h00000000; y17 = 32'h00000000; y16 = 32'h00000000; y15 = 32'h00000000; y14 = 32'h00000000;
	            y13 = 32'h00000000; y12 = 32'h00000000; y11 = 32'h00000000; y10 = 32'h00000000; y9 = 32'h00000000;  y8 = 32'h00000000;
		    y7 = 32'h00000000;  y6 = 32'h00000000;  y5 = 32'h00000000;  y4 = 32'h00000000;  y3 = 32'h00000000;  y2 = 32'h00000000;
		    y1 = 32'h00000000;  y0 = 32'h00000000;

		#10 y31 = 32'h00000000; y30 = 32'h00000000; y29 = 32'h00000000; y28 = 32'h00000000; y27 = 32'h00000000; y26 = 32'h00000000; 
	            y25 = 32'h00000000; y24 = 32'hFFFFFFFF; y23 = 32'h00000000; y22 = 32'h00000000; y21 = 32'h00000000; y20 = 32'h00000000;
		    y19 = 32'h00000000; y18 = 32'h00000000; y17 = 32'h00000000; y16 = 32'h00000000; y15 = 32'h00000000; y14 = 32'h00000000;
	            y13 = 32'h00000000; y12 = 32'h00000000; y11 = 32'h00000000; y10 = 32'h00000000; y9 = 32'h00000000;  y8 = 32'h00000000;
		    y7 = 32'h00000000;  y6 = 32'h00000000;  y5 = 32'h00000000;  y4 = 32'h00000000;  y3 = 32'h00000000;  y2 = 32'h00000000;
		    y1 = 32'h00000000;  y0 = 32'h00000000;


	//Select 11001
	#10 s4 = 1'b1; s3 = 1'b1; s2 = 1'b0; s1 = 1'b0; s0 = 1'b1;
		#10 y31 = 32'h00000000; y30 = 32'h00000000; y29 = 32'h00000000; y28 = 32'h00000000; y27 = 32'h00000000; y26 = 32'h00000000; 
	            y25 = 32'h00000000; y24 = 32'h00000000; y23 = 32'h00000000; y22 = 32'h00000000; y21 = 32'h00000000; y20 = 32'h00000000;
		    y19 = 32'h00000000; y18 = 32'h00000000; y17 = 32'h00000000; y16 = 32'h00000000; y15 = 32'h00000000; y14 = 32'h00000000;
	            y13 = 32'h00000000; y12 = 32'h00000000; y11 = 32'h00000000; y10 = 32'h00000000; y9 = 32'h00000000;  y8 = 32'h00000000;
		    y7 = 32'h00000000;  y6 = 32'h00000000;  y5 = 32'h00000000;  y4 = 32'h00000000;  y3 = 32'h00000000;  y2 = 32'h00000000;
		    y1 = 32'h00000000;  y0 = 32'h00000000;

		#10 y31 = 32'h00000000; y30 = 32'h00000000; y29 = 32'h00000000; y28 = 32'h00000000; y27 = 32'h00000000; y26 = 32'h00000000; 
	            y25 = 32'hFFFFFFFF; y24 = 32'h00000000; y23 = 32'h00000000; y22 = 32'h00000000; y21 = 32'h00000000; y20 = 32'h00000000;
		    y19 = 32'h00000000; y18 = 32'h00000000; y17 = 32'h00000000; y16 = 32'h00000000; y15 = 32'h00000000; y14 = 32'h00000000;
	            y13 = 32'h00000000; y12 = 32'h00000000; y11 = 32'h00000000; y10 = 32'h00000000; y9 = 32'h00000000;  y8 = 32'h00000000;
		    y7 = 32'h00000000;  y6 = 32'h00000000;  y5 = 32'h00000000;  y4 = 32'h00000000;  y3 = 32'h00000000;  y2 = 32'h00000000;
		    y1 = 32'h00000000;  y0 = 32'h00000000;

	//Select 11010
	#10 s4 = 1'b1; s3 = 1'b1; s2 = 1'b0; s1 = 1'b1; s0 = 1'b0;
		#10 y31 = 32'h00000000; y30 = 32'h00000000; y29 = 32'h00000000; y28 = 32'h00000000; y27 = 32'h00000000; y26 = 32'h00000000; 
	            y25 = 32'h00000000; y24 = 32'h00000000; y23 = 32'h00000000; y22 = 32'h00000000; y21 = 32'h00000000; y20 = 32'h00000000;
		    y19 = 32'h00000000; y18 = 32'h00000000; y17 = 32'h00000000; y16 = 32'h00000000; y15 = 32'h00000000; y14 = 32'h00000000;
	            y13 = 32'h00000000; y12 = 32'h00000000; y11 = 32'h00000000; y10 = 32'h00000000; y9 = 32'h00000000;  y8 = 32'h00000000;
		    y7 = 32'h00000000;  y6 = 32'h00000000;  y5 = 32'h00000000;  y4 = 32'h00000000;  y3 = 32'h00000000;  y2 = 32'h00000000;
		    y1 = 32'h00000000;  y0 = 32'h00000000;

		#10 y31 = 32'h00000000; y30 = 32'h00000000; y29 = 32'h00000000; y28 = 32'h00000000; y27 = 32'h00000000; y26 = 32'hFFFFFFFF; 
	            y25 = 32'h00000000; y24 = 32'h00000000; y23 = 32'h00000000; y22 = 32'h00000000; y21 = 32'h00000000; y20 = 32'h00000000;
		    y19 = 32'h00000000; y18 = 32'h00000000; y17 = 32'h00000000; y16 = 32'h00000000; y15 = 32'h00000000; y14 = 32'h00000000;
	            y13 = 32'h00000000; y12 = 32'h00000000; y11 = 32'h00000000; y10 = 32'h00000000; y9 = 32'h00000000;  y8 = 32'h00000000;
		    y7 = 32'h00000000;  y6 = 32'h00000000;  y5 = 32'h00000000;  y4 = 32'h00000000;  y3 = 32'h00000000;  y2 = 32'h00000000;
		    y1 = 32'h00000000;  y0 = 32'h00000000;

		

	//Select 11011
	#10 s4 = 1'b1; s3 = 1'b1; s2 = 1'b0; s1 = 1'b1; s0 = 1'b1;
		#10 y31 = 32'h00000000; y30 = 32'h00000000; y29 = 32'h00000000; y28 = 32'h00000000; y27 = 32'h00000000; y26 = 32'h00000000; 
	            y25 = 32'h00000000; y24 = 32'h00000000; y23 = 32'h00000000; y22 = 32'h00000000; y21 = 32'h00000000; y20 = 32'h00000000;
		    y19 = 32'h00000000; y18 = 32'h00000000; y17 = 32'h00000000; y16 = 32'h00000000; y15 = 32'h00000000; y14 = 32'h00000000;
	            y13 = 32'h00000000; y12 = 32'h00000000; y11 = 32'h00000000; y10 = 32'h00000000; y9 = 32'h00000000;  y8 = 32'h00000000;
		    y7 = 32'h00000000;  y6 = 32'h00000000;  y5 = 32'h00000000;  y4 = 32'h00000000;  y3 = 32'h00000000;  y2 = 32'h00000000;
		    y1 = 32'h00000000;  y0 = 32'h00000000;

		#10 y31 = 32'h00000000; y30 = 32'h00000000; y29 = 32'h00000000; y28 = 32'h00000000; y27 = 32'hFFFFFFFF; y26 = 32'h00000000; 
	            y25 = 32'h00000000; y24 = 32'h00000000; y23 = 32'h00000000; y22 = 32'h00000000; y21 = 32'h00000000; y20 = 32'h00000000;
		    y19 = 32'h00000000; y18 = 32'h00000000; y17 = 32'h00000000; y16 = 32'h00000000; y15 = 32'h00000000; y14 = 32'h00000000;
	            y13 = 32'h00000000; y12 = 32'h00000000; y11 = 32'h00000000; y10 = 32'h00000000; y9 = 32'h00000000;  y8 = 32'h00000000;
		    y7 = 32'h00000000;  y6 = 32'h00000000;  y5 = 32'h00000000;  y4 = 32'h00000000;  y3 = 32'h00000000;  y2 = 32'h00000000;
		    y1 = 32'h00000000;  y0 = 32'h00000000;

	//Select 11100
	#10 s4 = 1'b1; s3 = 1'b1; s2 = 1'b1; s1 = 1'b0; s0 = 1'b0;
		#10 y31 = 32'h00000000; y30 = 32'h00000000; y29 = 32'h00000000; y28 = 32'h00000000; y27 = 32'h00000000; y26 = 32'h00000000; 
	            y25 = 32'h00000000; y24 = 32'h00000000; y23 = 32'h00000000; y22 = 32'h00000000; y21 = 32'h00000000; y20 = 32'h00000000;
		    y19 = 32'h00000000; y18 = 32'h00000000; y17 = 32'h00000000; y16 = 32'h00000000; y15 = 32'h00000000; y14 = 32'h00000000;
	            y13 = 32'h00000000; y12 = 32'h00000000; y11 = 32'h00000000; y10 = 32'h00000000; y9 = 32'h00000000;  y8 = 32'h00000000;
		    y7 = 32'h00000000;  y6 = 32'h00000000;  y5 = 32'h00000000;  y4 = 32'h00000000;  y3 = 32'h00000000;  y2 = 32'h00000000;
		    y1 = 32'h00000000;  y0 = 32'h00000000;
	
		#10 y31 = 32'h00000000; y30 = 32'h00000000; y29 = 32'h00000000; y28 = 32'hFFFFFFFF; y27 = 32'h00000000; y26 = 32'h00000000; 
	            y25 = 32'h00000000; y24 = 32'h00000000; y23 = 32'h00000000; y22 = 32'h00000000; y21 = 32'h00000000; y20 = 32'h00000000;
		    y19 = 32'h00000000; y18 = 32'h00000000; y17 = 32'h00000000; y16 = 32'h00000000; y15 = 32'h00000000; y14 = 32'h00000000;
	            y13 = 32'h00000000; y12 = 32'h00000000; y11 = 32'h00000000; y10 = 32'h00000000; y9 = 32'h00000000;  y8 = 32'h00000000;
		    y7 = 32'h00000000;  y6 = 32'h00000000;  y5 = 32'h00000000;  y4 = 32'h00000000;  y3 = 32'h00000000;  y2 = 32'h00000000;
		    y1 = 32'h00000000;  y0 = 32'h00000000;

	//Select 11101
	#10 s4 = 1'b1; s3 = 1'b1; s2 = 1'b1; s1 = 1'b0; s0 = 1'b1;
		#10 y31 = 32'h00000000; y30 = 32'h00000000; y29 = 32'h00000000; y28 = 32'h00000000; y27 = 32'h00000000; y26 = 32'h00000000; 
	            y25 = 32'h00000000; y24 = 32'h00000000; y23 = 32'h00000000; y22 = 32'h00000000; y21 = 32'h00000000; y20 = 32'h00000000;
		    y19 = 32'h00000000; y18 = 32'h00000000; y17 = 32'h00000000; y16 = 32'h00000000; y15 = 32'h00000000; y14 = 32'h00000000;
	            y13 = 32'h00000000; y12 = 32'h00000000; y11 = 32'h00000000; y10 = 32'h00000000; y9 = 32'h00000000;  y8 = 32'h00000000;
		    y7 = 32'h00000000;  y6 = 32'h00000000;  y5 = 32'h00000000;  y4 = 32'h00000000;  y3 = 32'h00000000;  y2 = 32'h00000000;
		    y1 = 32'h00000000;  y0 = 32'h00000000;

		#10 y31 = 32'h00000000; y30 = 32'h00000000; y29 = 32'hFFFFFFFF; y28 = 32'h00000000; y27 = 32'h00000000; y26 = 32'h00000000; 
	            y25 = 32'h00000000; y24 = 32'h00000000; y23 = 32'h00000000; y22 = 32'h00000000; y21 = 32'h00000000; y20 = 32'h00000000;
		    y19 = 32'h00000000; y18 = 32'h00000000; y17 = 32'h00000000; y16 = 32'h00000000; y15 = 32'h00000000; y14 = 32'h00000000;
	            y13 = 32'h00000000; y12 = 32'h00000000; y11 = 32'h00000000; y10 = 32'h00000000; y9 = 32'h00000000;  y8 = 32'h00000000;
		    y7 = 32'h00000000;  y6 = 32'h00000000;  y5 = 32'h00000000;  y4 = 32'h00000000;  y3 = 32'h00000000;  y2 = 32'h00000000;
		    y1 = 32'h00000000;  y0 = 32'h00000000;

	//Select 11110
	#10 s4 = 1'b1; s3 = 1'b1; s2 = 1'b1; s1 = 1'b1; s0 = 1'b0;
		#10 y31 = 32'h00000000; y30 = 32'h00000000; y29 = 32'h00000000; y28 = 32'h00000000; y27 = 32'h00000000; y26 = 32'h00000000; 
	            y25 = 32'h00000000; y24 = 32'h00000000; y23 = 32'h00000000; y22 = 32'h00000000; y21 = 32'h00000000; y20 = 32'h00000000;
		    y19 = 32'h00000000; y18 = 32'h00000000; y17 = 32'h00000000; y16 = 32'h00000000; y15 = 32'h00000000; y14 = 32'h00000000;
	            y13 = 32'h00000000; y12 = 32'h00000000; y11 = 32'h00000000; y10 = 32'h00000000; y9 = 32'h00000000;  y8 = 32'h00000000;
		    y7 = 32'h00000000;  y6 = 32'h00000000;  y5 = 32'h00000000;  y4 = 32'h00000000;  y3 = 32'h00000000;  y2 = 32'h00000000;
		    y1 = 32'h00000000;  y0 = 32'h00000000;

		#10 y31 = 32'h00000000; y30 = 32'hFFFFFFFF; y29 = 32'h00000000; y28 = 32'h00000000; y27 = 32'h00000000; y26 = 32'h00000000; 
	            y25 = 32'h00000000; y24 = 32'h00000000; y23 = 32'h00000000; y22 = 32'h00000000; y21 = 32'h00000000; y20 = 32'h00000000;
		    y19 = 32'h00000000; y18 = 32'h00000000; y17 = 32'h00000000; y16 = 32'h00000000; y15 = 32'h00000000; y14 = 32'h00000000;
	            y13 = 32'h00000000; y12 = 32'h00000000; y11 = 32'h00000000; y10 = 32'h00000000; y9 = 32'h00000000;  y8 = 32'h00000000;
		    y7 = 32'h00000000;  y6 = 32'h00000000;  y5 = 32'h00000000;  y4 = 32'h00000000;  y3 = 32'h00000000;  y2 = 32'h00000000;
		    y1 = 32'h00000000;  y0 = 32'h00000000;

	//Select 11111
	#10 s4 = 1'b1; s3 = 1'b1; s2 = 1'b1; s1 = 1'b0; s0 = 1'b1;
		#10 y31 = 32'h00000000; y30 = 32'h00000000; y29 = 32'h00000000; y28 = 32'h00000000; y27 = 32'h00000000; y26 = 32'h00000000; 
	            y25 = 32'h00000000; y24 = 32'h00000000; y23 = 32'h00000000; y22 = 32'h00000000; y21 = 32'h00000000; y20 = 32'h00000000;
		    y19 = 32'h00000000; y18 = 32'h00000000; y17 = 32'h00000000; y16 = 32'h00000000; y15 = 32'h00000000; y14 = 32'h00000000;
	            y13 = 32'h00000000; y12 = 32'h00000000; y11 = 32'h00000000; y10 = 32'h00000000; y9 = 32'h00000000;  y8 = 32'h00000000;
		    y7 = 32'h00000000;  y6 = 32'h00000000;  y5 = 32'h00000000;  y4 = 32'h00000000;  y3 = 32'h00000000;  y2 = 32'h00000000;
		    y1 = 32'h00000000;  y0 = 32'h00000000;

		#10 y31 = 32'hFFFFFFFF; y30 = 32'h00000000; y29 = 32'h00000000; y28 = 32'h00000000; y27 = 32'h00000000; y26 = 32'h00000000; 
	            y25 = 32'h00000000; y24 = 32'h00000000; y23 = 32'h00000000; y22 = 32'h00000000; y21 = 32'h00000000; y20 = 32'h00000000;
		    y19 = 32'h00000000; y18 = 32'h00000000; y17 = 32'h00000000; y16 = 32'h00000000; y15 = 32'h00000000; y14 = 32'h00000000;
	            y13 = 32'h00000000; y12 = 32'h00000000; y11 = 32'h00000000; y10 = 32'h00000000; y9 = 32'h00000000;  y8 = 32'h00000000;
		    y7 = 32'h00000000;  y6 = 32'h00000000;  y5 = 32'h00000000;  y4 = 32'h00000000;  y3 = 32'h00000000;  y2 = 32'h00000000;
		    y1 = 32'h00000000;  y0 = 32'h00000000;

	#10 $stop;
  end


initial
  begin
	$display("		  time 		y31 y30 y29 y28 y27 y26 y25 y24 y23" + 
			" y22 y21 y20 y19 y18 y17 y16 y15 y14 y13 y12 y11 y10 y9 y8 y7 " +
			"y6 y5 y4 y3 y2 y1 y0 s4 s3 s2 s1 s0 		z");
	$monitor($time,, y31,, y30,, y29,, y28,, y27,, y26,, y25,, y24,, y23,, y22,, y21,, y20,, y19,, 
			y18,, y17,, y16,, y15,, y14,, y13,, y12,, y11,, y10,, y9,, y8,, y7,, y6,, y5,, 
			y4,, y3,, y2,, y1,, y0,, s4,, s3,, s2,, s1,, s0,,,,,, z);
  end

endmodule